magic
tech scmos
timestamp 1593933729
<< nsubstratencontact >>
rect -130 35 -122 47
rect 59 4 67 16
<< rnwell >>
rect -122 35 67 47
rect 55 31 67 35
rect -130 19 67 31
rect -130 16 -118 19
rect -130 4 59 16
<< pseudo_nwr >>
rect -131 47 68 48
rect -131 35 -130 47
rect -131 31 55 35
rect -131 4 -130 31
rect 67 19 68 47
rect -118 16 68 19
rect 67 4 68 16
rect -131 -72 68 4
<< labels >>
rlabel nsubstratencontact 64 13 64 13 7 b
rlabel nsubstratencontact -127 43 -127 43 4 a
<< end >>
