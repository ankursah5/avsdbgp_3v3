* SPICE3 file created from bgr1.ext - technology: scmos

.option scale=0.1u

Q1000 0 0 N006 PNP
Q1001 0 0 vctat PNP
Q1002 0 0 N007 PNP
Q1003 0 0 N007 PNP
Q1004 0 0 N007 PNP
Q1005 0 0 N007 PNP
Q1006 0 0 N007 PNP
Q1007 0 0 N007 PNP
Q1008 0 0 N007 PNP
Q1009 0 0 N007 PNP
M1010 N001 N002 N002 N001 pfet w=100 l=50
+  ad=6000 pd=720 as=2000 ps=240
Q1011 0 N001 N001 PNP
M1012 0 N003 N004 0 nfet w=200 l=50
+  ad=21340 pd=4330 as=4144 ps=488
M1013 N003 N003 N006 0 nfet w=100 l=50
+  ad=2000 pd=240 as=2000 ps=240
M1014 N005 N003 N002 0 nfet w=100 l=50
+  ad=2120 pd=284 as=2300 ps=310
M1015 N002 N004 0 0 nfet w=20 l=20
+  ad=0 pd=0 as=0 ps=0
R0 N005 N007 nwellResistor w=12 l=103
Q1016 0 N001 vref PNP
M1017 N001 N002 vref N001 pfet w=100 l=50
+  ad=0 pd=0 as=2000 ps=240
R1 N001 N004 nwellResistor w=12 l=15428
R2 vref vctat nwellResistor w=12 l=1275
Q1018 0 N001 N002 PNP
M1019 N003 N002 N001 N001 pfet w=100 l=50
+  ad=2000 pd=240 as=0 ps=0
C0 N002 N001 7.36fF
C1 a_221_n129# 0 12.07fF **FLOATING
C2 N004 0 2.57fF
C3 N003 0 8.80fF
C4 a_n999_n265# 0 143.33fF **FLOATING
C5 N001 0 61.60fF
C6 N007 0 12.42fF
